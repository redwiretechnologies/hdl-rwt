// Tags are 7-bits wide.
localparam RWT_TAG_TIME = 7'd01;
localparam RWT_TAG_PPS = 7'd02;
localparam RWT_TAG_OVERFLOW = 7'd03;

localparam RWT_TAG_HOLD = 7'd04;
localparam RWT_TAG_SOB = 7'd05;
localparam RWT_TAG_EOB = 7'd06;
