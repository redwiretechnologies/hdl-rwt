// SPDX-License-Identifier: Apache-2.0

`ifndef RWT_SV
`define RWT_SV

`include "rwt_parse_utils.sv"
`include "rwt_axis.sv"
`include "rwt_axi4lite_lib.sv"
`include "rwt_axis_tag_pkt.sv"
`include "rwt_up_lib.sv"
`include "rwt_adc_lib.sv"
`include "rwt_dac_lib.sv"

`endif
