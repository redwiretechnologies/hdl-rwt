// Tags are 7-bits wide.
localparam RWT_TAG_TIME = 'd01;
localparam RWT_TAG_PPS = 'd02;
localparam RWT_TAG_OVERFLOW = 'd03;

localparam RWT_TAG_HOLD = 'd04;
localparam RWT_TAG_SOB = 'd05;
localparam RWT_TAG_EOB = 'd06;
